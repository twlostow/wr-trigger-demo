library ieee;
use ieee.std_logic_1164.all;
package pack_unpack_pkg is
procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic);
procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector);
end pack_unpack_pkg;
package body pack_unpack_pkg is
procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
end f_unpack2;

procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
end f_unpack2;

procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
end f_unpack2;

procedure f_unpack2 (
x: in std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
end f_unpack2;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
end f_unpack3;

procedure f_unpack3 (
x: in std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
end f_unpack3;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
end f_unpack4;

procedure f_unpack4 (
x: in std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
end f_unpack4;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
end f_unpack5;

procedure f_unpack5 (
x: in std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
end f_unpack5;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
q5 :=x(0+1+1+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
q5 :=x(0+q0'length+1+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
q5 :=x(0+1+q1'length+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
q5 :=x(0+q0'length+q1'length+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
q5 :=x(0+1+1+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
q5 :=x(0+q0'length+1+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
q5 :=x(0+1+q1'length+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
q5 :=x(0+q0'length+q1'length+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
q5 :=x(0+1+1+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
q5 :=x(0+q0'length+1+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
q5 :=x(0+1+q1'length+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
q5 :=x(0+q0'length+q1'length+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
q5 :=x(0+1+1+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
q5 :=x(0+q0'length+1+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
q5 :=x(0+1+q1'length+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(0+q0'length+q1'length+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
q5 :=x(0+1+1+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
q5 :=x(0+q0'length+1+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
q5 :=x(0+1+q1'length+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
q5 :=x(0+q0'length+q1'length+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
q5 :=x(0+1+1+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
q5 :=x(0+q0'length+1+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
q5 :=x(0+1+q1'length+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
q5 :=x(0+q0'length+q1'length+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
q5 :=x(0+1+1+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
q5 :=x(0+q0'length+1+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
q5 :=x(0+1+q1'length+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
q5 :=x(0+q0'length+q1'length+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
q5 :=x(0+1+1+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
q5 :=x(0+q0'length+1+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
q5 :=x(0+1+q1'length+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(0+q0'length+q1'length+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
q5 :=x(-1+1+1+1+1+1+q5'length downto 0+1+1+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
q5 :=x(-1+q0'length+1+1+1+1+q5'length downto 0+q0'length+1+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
q5 :=x(-1+1+q1'length+1+1+1+q5'length downto 0+1+q1'length+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
q5 :=x(-1+q0'length+q1'length+1+1+1+q5'length downto 0+q0'length+q1'length+1+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
q5 :=x(-1+1+1+q2'length+1+1+q5'length downto 0+1+1+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
q5 :=x(-1+q0'length+1+q2'length+1+1+q5'length downto 0+q0'length+1+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
q5 :=x(-1+1+q1'length+q2'length+1+1+q5'length downto 0+1+q1'length+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
q5 :=x(-1+q0'length+q1'length+q2'length+1+1+q5'length downto 0+q0'length+q1'length+q2'length+1+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
q5 :=x(-1+1+1+1+q3'length+1+q5'length downto 0+1+1+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
q5 :=x(-1+q0'length+1+1+q3'length+1+q5'length downto 0+q0'length+1+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
q5 :=x(-1+1+q1'length+1+q3'length+1+q5'length downto 0+1+q1'length+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
q5 :=x(-1+q0'length+q1'length+1+q3'length+1+q5'length downto 0+q0'length+q1'length+1+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
q5 :=x(-1+1+1+q2'length+q3'length+1+q5'length downto 0+1+1+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
q5 :=x(-1+q0'length+1+q2'length+q3'length+1+q5'length downto 0+q0'length+1+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
q5 :=x(-1+1+q1'length+q2'length+q3'length+1+q5'length downto 0+1+q1'length+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(-1+q0'length+q1'length+q2'length+q3'length+1+q5'length downto 0+q0'length+q1'length+q2'length+q3'length+1);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
q5 :=x(-1+1+1+1+1+q4'length+q5'length downto 0+1+1+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
q5 :=x(-1+q0'length+1+1+1+q4'length+q5'length downto 0+q0'length+1+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
q5 :=x(-1+1+q1'length+1+1+q4'length+q5'length downto 0+1+q1'length+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
q5 :=x(-1+q0'length+q1'length+1+1+q4'length+q5'length downto 0+q0'length+q1'length+1+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
q5 :=x(-1+1+1+q2'length+1+q4'length+q5'length downto 0+1+1+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
q5 :=x(-1+q0'length+1+q2'length+1+q4'length+q5'length downto 0+q0'length+1+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
q5 :=x(-1+1+q1'length+q2'length+1+q4'length+q5'length downto 0+1+q1'length+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
q5 :=x(-1+q0'length+q1'length+q2'length+1+q4'length+q5'length downto 0+q0'length+q1'length+q2'length+1+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
q5 :=x(-1+1+1+1+q3'length+q4'length+q5'length downto 0+1+1+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
q5 :=x(-1+q0'length+1+1+q3'length+q4'length+q5'length downto 0+q0'length+1+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
q5 :=x(-1+1+q1'length+1+q3'length+q4'length+q5'length downto 0+1+q1'length+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
q5 :=x(-1+q0'length+q1'length+1+q3'length+q4'length+q5'length downto 0+q0'length+q1'length+1+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
q5 :=x(-1+1+1+q2'length+q3'length+q4'length+q5'length downto 0+1+1+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
q5 :=x(-1+q0'length+1+q2'length+q3'length+q4'length+q5'length downto 0+q0'length+1+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
q5 :=x(-1+1+q1'length+q2'length+q3'length+q4'length+q5'length downto 0+1+q1'length+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack6 (
x: in std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length+q5'length downto 0+q0'length+q1'length+q2'length+q3'length+q4'length);
end f_unpack6;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
q5 :=x(0+1+1+1+1+1);
q6 :=x(0+1+1+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
q5 :=x(0+q0'length+1+1+1+1);
q6 :=x(0+q0'length+1+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
q5 :=x(0+1+q1'length+1+1+1);
q6 :=x(0+1+q1'length+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
q5 :=x(0+q0'length+q1'length+1+1+1);
q6 :=x(0+q0'length+q1'length+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
q5 :=x(0+1+1+q2'length+1+1);
q6 :=x(0+1+1+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
q5 :=x(0+q0'length+1+q2'length+1+1);
q6 :=x(0+q0'length+1+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
q5 :=x(0+1+q1'length+q2'length+1+1);
q6 :=x(0+1+q1'length+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
q5 :=x(0+q0'length+q1'length+q2'length+1+1);
q6 :=x(0+q0'length+q1'length+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
q5 :=x(0+1+1+1+q3'length+1);
q6 :=x(0+1+1+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
q5 :=x(0+q0'length+1+1+q3'length+1);
q6 :=x(0+q0'length+1+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
q5 :=x(0+1+q1'length+1+q3'length+1);
q6 :=x(0+1+q1'length+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
q5 :=x(0+q0'length+q1'length+1+q3'length+1);
q6 :=x(0+q0'length+q1'length+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
q5 :=x(0+1+1+q2'length+q3'length+1);
q6 :=x(0+1+1+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
q5 :=x(0+q0'length+1+q2'length+q3'length+1);
q6 :=x(0+q0'length+1+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
q5 :=x(0+1+q1'length+q2'length+q3'length+1);
q6 :=x(0+1+q1'length+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(0+q0'length+q1'length+q2'length+q3'length+1);
q6 :=x(0+q0'length+q1'length+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
q5 :=x(0+1+1+1+1+q4'length);
q6 :=x(0+1+1+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
q5 :=x(0+q0'length+1+1+1+q4'length);
q6 :=x(0+q0'length+1+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
q5 :=x(0+1+q1'length+1+1+q4'length);
q6 :=x(0+1+q1'length+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
q5 :=x(0+q0'length+q1'length+1+1+q4'length);
q6 :=x(0+q0'length+q1'length+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
q5 :=x(0+1+1+q2'length+1+q4'length);
q6 :=x(0+1+1+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
q5 :=x(0+q0'length+1+q2'length+1+q4'length);
q6 :=x(0+q0'length+1+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
q5 :=x(0+1+q1'length+q2'length+1+q4'length);
q6 :=x(0+1+q1'length+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
q5 :=x(0+q0'length+q1'length+q2'length+1+q4'length);
q6 :=x(0+q0'length+q1'length+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
q5 :=x(0+1+1+1+q3'length+q4'length);
q6 :=x(0+1+1+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
q5 :=x(0+q0'length+1+1+q3'length+q4'length);
q6 :=x(0+q0'length+1+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
q5 :=x(0+1+q1'length+1+q3'length+q4'length);
q6 :=x(0+1+q1'length+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
q5 :=x(0+q0'length+q1'length+1+q3'length+q4'length);
q6 :=x(0+q0'length+q1'length+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
q5 :=x(0+1+1+q2'length+q3'length+q4'length);
q6 :=x(0+1+1+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
q5 :=x(0+q0'length+1+q2'length+q3'length+q4'length);
q6 :=x(0+q0'length+1+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
q5 :=x(0+1+q1'length+q2'length+q3'length+q4'length);
q6 :=x(0+1+q1'length+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(0+q0'length+q1'length+q2'length+q3'length+q4'length);
q6 :=x(0+q0'length+q1'length+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
q5 :=x(-1+1+1+1+1+1+q5'length downto 0+1+1+1+1+1);
q6 :=x(0+1+1+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
q5 :=x(-1+q0'length+1+1+1+1+q5'length downto 0+q0'length+1+1+1+1);
q6 :=x(0+q0'length+1+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
q5 :=x(-1+1+q1'length+1+1+1+q5'length downto 0+1+q1'length+1+1+1);
q6 :=x(0+1+q1'length+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
q5 :=x(-1+q0'length+q1'length+1+1+1+q5'length downto 0+q0'length+q1'length+1+1+1);
q6 :=x(0+q0'length+q1'length+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
q5 :=x(-1+1+1+q2'length+1+1+q5'length downto 0+1+1+q2'length+1+1);
q6 :=x(0+1+1+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
q5 :=x(-1+q0'length+1+q2'length+1+1+q5'length downto 0+q0'length+1+q2'length+1+1);
q6 :=x(0+q0'length+1+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
q5 :=x(-1+1+q1'length+q2'length+1+1+q5'length downto 0+1+q1'length+q2'length+1+1);
q6 :=x(0+1+q1'length+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
q5 :=x(-1+q0'length+q1'length+q2'length+1+1+q5'length downto 0+q0'length+q1'length+q2'length+1+1);
q6 :=x(0+q0'length+q1'length+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
q5 :=x(-1+1+1+1+q3'length+1+q5'length downto 0+1+1+1+q3'length+1);
q6 :=x(0+1+1+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
q5 :=x(-1+q0'length+1+1+q3'length+1+q5'length downto 0+q0'length+1+1+q3'length+1);
q6 :=x(0+q0'length+1+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
q5 :=x(-1+1+q1'length+1+q3'length+1+q5'length downto 0+1+q1'length+1+q3'length+1);
q6 :=x(0+1+q1'length+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
q5 :=x(-1+q0'length+q1'length+1+q3'length+1+q5'length downto 0+q0'length+q1'length+1+q3'length+1);
q6 :=x(0+q0'length+q1'length+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
q5 :=x(-1+1+1+q2'length+q3'length+1+q5'length downto 0+1+1+q2'length+q3'length+1);
q6 :=x(0+1+1+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
q5 :=x(-1+q0'length+1+q2'length+q3'length+1+q5'length downto 0+q0'length+1+q2'length+q3'length+1);
q6 :=x(0+q0'length+1+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
q5 :=x(-1+1+q1'length+q2'length+q3'length+1+q5'length downto 0+1+q1'length+q2'length+q3'length+1);
q6 :=x(0+1+q1'length+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(-1+q0'length+q1'length+q2'length+q3'length+1+q5'length downto 0+q0'length+q1'length+q2'length+q3'length+1);
q6 :=x(0+q0'length+q1'length+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
q5 :=x(-1+1+1+1+1+q4'length+q5'length downto 0+1+1+1+1+q4'length);
q6 :=x(0+1+1+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
q5 :=x(-1+q0'length+1+1+1+q4'length+q5'length downto 0+q0'length+1+1+1+q4'length);
q6 :=x(0+q0'length+1+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
q5 :=x(-1+1+q1'length+1+1+q4'length+q5'length downto 0+1+q1'length+1+1+q4'length);
q6 :=x(0+1+q1'length+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
q5 :=x(-1+q0'length+q1'length+1+1+q4'length+q5'length downto 0+q0'length+q1'length+1+1+q4'length);
q6 :=x(0+q0'length+q1'length+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
q5 :=x(-1+1+1+q2'length+1+q4'length+q5'length downto 0+1+1+q2'length+1+q4'length);
q6 :=x(0+1+1+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
q5 :=x(-1+q0'length+1+q2'length+1+q4'length+q5'length downto 0+q0'length+1+q2'length+1+q4'length);
q6 :=x(0+q0'length+1+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
q5 :=x(-1+1+q1'length+q2'length+1+q4'length+q5'length downto 0+1+q1'length+q2'length+1+q4'length);
q6 :=x(0+1+q1'length+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
q5 :=x(-1+q0'length+q1'length+q2'length+1+q4'length+q5'length downto 0+q0'length+q1'length+q2'length+1+q4'length);
q6 :=x(0+q0'length+q1'length+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
q5 :=x(-1+1+1+1+q3'length+q4'length+q5'length downto 0+1+1+1+q3'length+q4'length);
q6 :=x(0+1+1+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
q5 :=x(-1+q0'length+1+1+q3'length+q4'length+q5'length downto 0+q0'length+1+1+q3'length+q4'length);
q6 :=x(0+q0'length+1+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
q5 :=x(-1+1+q1'length+1+q3'length+q4'length+q5'length downto 0+1+q1'length+1+q3'length+q4'length);
q6 :=x(0+1+q1'length+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
q5 :=x(-1+q0'length+q1'length+1+q3'length+q4'length+q5'length downto 0+q0'length+q1'length+1+q3'length+q4'length);
q6 :=x(0+q0'length+q1'length+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
q5 :=x(-1+1+1+q2'length+q3'length+q4'length+q5'length downto 0+1+1+q2'length+q3'length+q4'length);
q6 :=x(0+1+1+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
q5 :=x(-1+q0'length+1+q2'length+q3'length+q4'length+q5'length downto 0+q0'length+1+q2'length+q3'length+q4'length);
q6 :=x(0+q0'length+1+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
q5 :=x(-1+1+q1'length+q2'length+q3'length+q4'length+q5'length downto 0+1+q1'length+q2'length+q3'length+q4'length);
q6 :=x(0+1+q1'length+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length+q5'length downto 0+q0'length+q1'length+q2'length+q3'length+q4'length);
q6 :=x(0+q0'length+q1'length+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
q5 :=x(0+1+1+1+1+1);
q6 :=x(-1+1+1+1+1+1+1+q6'length downto 0+1+1+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
q5 :=x(0+q0'length+1+1+1+1);
q6 :=x(-1+q0'length+1+1+1+1+1+q6'length downto 0+q0'length+1+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
q5 :=x(0+1+q1'length+1+1+1);
q6 :=x(-1+1+q1'length+1+1+1+1+q6'length downto 0+1+q1'length+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
q5 :=x(0+q0'length+q1'length+1+1+1);
q6 :=x(-1+q0'length+q1'length+1+1+1+1+q6'length downto 0+q0'length+q1'length+1+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
q5 :=x(0+1+1+q2'length+1+1);
q6 :=x(-1+1+1+q2'length+1+1+1+q6'length downto 0+1+1+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
q5 :=x(0+q0'length+1+q2'length+1+1);
q6 :=x(-1+q0'length+1+q2'length+1+1+1+q6'length downto 0+q0'length+1+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
q5 :=x(0+1+q1'length+q2'length+1+1);
q6 :=x(-1+1+q1'length+q2'length+1+1+1+q6'length downto 0+1+q1'length+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
q5 :=x(0+q0'length+q1'length+q2'length+1+1);
q6 :=x(-1+q0'length+q1'length+q2'length+1+1+1+q6'length downto 0+q0'length+q1'length+q2'length+1+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
q5 :=x(0+1+1+1+q3'length+1);
q6 :=x(-1+1+1+1+q3'length+1+1+q6'length downto 0+1+1+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
q5 :=x(0+q0'length+1+1+q3'length+1);
q6 :=x(-1+q0'length+1+1+q3'length+1+1+q6'length downto 0+q0'length+1+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
q5 :=x(0+1+q1'length+1+q3'length+1);
q6 :=x(-1+1+q1'length+1+q3'length+1+1+q6'length downto 0+1+q1'length+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
q5 :=x(0+q0'length+q1'length+1+q3'length+1);
q6 :=x(-1+q0'length+q1'length+1+q3'length+1+1+q6'length downto 0+q0'length+q1'length+1+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
q5 :=x(0+1+1+q2'length+q3'length+1);
q6 :=x(-1+1+1+q2'length+q3'length+1+1+q6'length downto 0+1+1+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
q5 :=x(0+q0'length+1+q2'length+q3'length+1);
q6 :=x(-1+q0'length+1+q2'length+q3'length+1+1+q6'length downto 0+q0'length+1+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
q5 :=x(0+1+q1'length+q2'length+q3'length+1);
q6 :=x(-1+1+q1'length+q2'length+q3'length+1+1+q6'length downto 0+1+q1'length+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(0+q0'length+q1'length+q2'length+q3'length+1);
q6 :=x(-1+q0'length+q1'length+q2'length+q3'length+1+1+q6'length downto 0+q0'length+q1'length+q2'length+q3'length+1+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
q5 :=x(0+1+1+1+1+q4'length);
q6 :=x(-1+1+1+1+1+q4'length+1+q6'length downto 0+1+1+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
q5 :=x(0+q0'length+1+1+1+q4'length);
q6 :=x(-1+q0'length+1+1+1+q4'length+1+q6'length downto 0+q0'length+1+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
q5 :=x(0+1+q1'length+1+1+q4'length);
q6 :=x(-1+1+q1'length+1+1+q4'length+1+q6'length downto 0+1+q1'length+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
q5 :=x(0+q0'length+q1'length+1+1+q4'length);
q6 :=x(-1+q0'length+q1'length+1+1+q4'length+1+q6'length downto 0+q0'length+q1'length+1+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
q5 :=x(0+1+1+q2'length+1+q4'length);
q6 :=x(-1+1+1+q2'length+1+q4'length+1+q6'length downto 0+1+1+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
q5 :=x(0+q0'length+1+q2'length+1+q4'length);
q6 :=x(-1+q0'length+1+q2'length+1+q4'length+1+q6'length downto 0+q0'length+1+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
q5 :=x(0+1+q1'length+q2'length+1+q4'length);
q6 :=x(-1+1+q1'length+q2'length+1+q4'length+1+q6'length downto 0+1+q1'length+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
q5 :=x(0+q0'length+q1'length+q2'length+1+q4'length);
q6 :=x(-1+q0'length+q1'length+q2'length+1+q4'length+1+q6'length downto 0+q0'length+q1'length+q2'length+1+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
q5 :=x(0+1+1+1+q3'length+q4'length);
q6 :=x(-1+1+1+1+q3'length+q4'length+1+q6'length downto 0+1+1+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
q5 :=x(0+q0'length+1+1+q3'length+q4'length);
q6 :=x(-1+q0'length+1+1+q3'length+q4'length+1+q6'length downto 0+q0'length+1+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
q5 :=x(0+1+q1'length+1+q3'length+q4'length);
q6 :=x(-1+1+q1'length+1+q3'length+q4'length+1+q6'length downto 0+1+q1'length+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
q5 :=x(0+q0'length+q1'length+1+q3'length+q4'length);
q6 :=x(-1+q0'length+q1'length+1+q3'length+q4'length+1+q6'length downto 0+q0'length+q1'length+1+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
q5 :=x(0+1+1+q2'length+q3'length+q4'length);
q6 :=x(-1+1+1+q2'length+q3'length+q4'length+1+q6'length downto 0+1+1+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
q5 :=x(0+q0'length+1+q2'length+q3'length+q4'length);
q6 :=x(-1+q0'length+1+q2'length+q3'length+q4'length+1+q6'length downto 0+q0'length+1+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
q5 :=x(0+1+q1'length+q2'length+q3'length+q4'length);
q6 :=x(-1+1+q1'length+q2'length+q3'length+q4'length+1+q6'length downto 0+1+q1'length+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(0+q0'length+q1'length+q2'length+q3'length+q4'length);
q6 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length+1+q6'length downto 0+q0'length+q1'length+q2'length+q3'length+q4'length+1);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(0+1+1+1+1);
q5 :=x(-1+1+1+1+1+1+q5'length downto 0+1+1+1+1+1);
q6 :=x(-1+1+1+1+1+1+q5'length+q6'length downto 0+1+1+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+1);
q5 :=x(-1+q0'length+1+1+1+1+q5'length downto 0+q0'length+1+1+1+1);
q6 :=x(-1+q0'length+1+1+1+1+q5'length+q6'length downto 0+q0'length+1+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+1);
q5 :=x(-1+1+q1'length+1+1+1+q5'length downto 0+1+q1'length+1+1+1);
q6 :=x(-1+1+q1'length+1+1+1+q5'length+q6'length downto 0+1+q1'length+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+1);
q5 :=x(-1+q0'length+q1'length+1+1+1+q5'length downto 0+q0'length+q1'length+1+1+1);
q6 :=x(-1+q0'length+q1'length+1+1+1+q5'length+q6'length downto 0+q0'length+q1'length+1+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+1);
q5 :=x(-1+1+1+q2'length+1+1+q5'length downto 0+1+1+q2'length+1+1);
q6 :=x(-1+1+1+q2'length+1+1+q5'length+q6'length downto 0+1+1+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+1);
q5 :=x(-1+q0'length+1+q2'length+1+1+q5'length downto 0+q0'length+1+q2'length+1+1);
q6 :=x(-1+q0'length+1+q2'length+1+1+q5'length+q6'length downto 0+q0'length+1+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+1);
q5 :=x(-1+1+q1'length+q2'length+1+1+q5'length downto 0+1+q1'length+q2'length+1+1);
q6 :=x(-1+1+q1'length+q2'length+1+1+q5'length+q6'length downto 0+1+q1'length+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+1);
q5 :=x(-1+q0'length+q1'length+q2'length+1+1+q5'length downto 0+q0'length+q1'length+q2'length+1+1);
q6 :=x(-1+q0'length+q1'length+q2'length+1+1+q5'length+q6'length downto 0+q0'length+q1'length+q2'length+1+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(0+1+1+1+q3'length);
q5 :=x(-1+1+1+1+q3'length+1+q5'length downto 0+1+1+1+q3'length+1);
q6 :=x(-1+1+1+1+q3'length+1+q5'length+q6'length downto 0+1+1+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(0+q0'length+1+1+q3'length);
q5 :=x(-1+q0'length+1+1+q3'length+1+q5'length downto 0+q0'length+1+1+q3'length+1);
q6 :=x(-1+q0'length+1+1+q3'length+1+q5'length+q6'length downto 0+q0'length+1+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(0+1+q1'length+1+q3'length);
q5 :=x(-1+1+q1'length+1+q3'length+1+q5'length downto 0+1+q1'length+1+q3'length+1);
q6 :=x(-1+1+q1'length+1+q3'length+1+q5'length+q6'length downto 0+1+q1'length+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(0+q0'length+q1'length+1+q3'length);
q5 :=x(-1+q0'length+q1'length+1+q3'length+1+q5'length downto 0+q0'length+q1'length+1+q3'length+1);
q6 :=x(-1+q0'length+q1'length+1+q3'length+1+q5'length+q6'length downto 0+q0'length+q1'length+1+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(0+1+1+q2'length+q3'length);
q5 :=x(-1+1+1+q2'length+q3'length+1+q5'length downto 0+1+1+q2'length+q3'length+1);
q6 :=x(-1+1+1+q2'length+q3'length+1+q5'length+q6'length downto 0+1+1+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(0+q0'length+1+q2'length+q3'length);
q5 :=x(-1+q0'length+1+q2'length+q3'length+1+q5'length downto 0+q0'length+1+q2'length+q3'length+1);
q6 :=x(-1+q0'length+1+q2'length+q3'length+1+q5'length+q6'length downto 0+q0'length+1+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(0+1+q1'length+q2'length+q3'length);
q5 :=x(-1+1+q1'length+q2'length+q3'length+1+q5'length downto 0+1+q1'length+q2'length+q3'length+1);
q6 :=x(-1+1+q1'length+q2'length+q3'length+1+q5'length+q6'length downto 0+1+q1'length+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(-1+q0'length+q1'length+q2'length+q3'length+1+q5'length downto 0+q0'length+q1'length+q2'length+q3'length+1);
q6 :=x(-1+q0'length+q1'length+q2'length+q3'length+1+q5'length+q6'length downto 0+q0'length+q1'length+q2'length+q3'length+1+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(0+1+1+1);
q4 :=x(-1+1+1+1+1+q4'length downto 0+1+1+1+1);
q5 :=x(-1+1+1+1+1+q4'length+q5'length downto 0+1+1+1+1+q4'length);
q6 :=x(-1+1+1+1+1+q4'length+q5'length+q6'length downto 0+1+1+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+1+q4'length downto 0+q0'length+1+1+1);
q5 :=x(-1+q0'length+1+1+1+q4'length+q5'length downto 0+q0'length+1+1+1+q4'length);
q6 :=x(-1+q0'length+1+1+1+q4'length+q5'length+q6'length downto 0+q0'length+1+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+1+q4'length downto 0+1+q1'length+1+1);
q5 :=x(-1+1+q1'length+1+1+q4'length+q5'length downto 0+1+q1'length+1+1+q4'length);
q6 :=x(-1+1+q1'length+1+1+q4'length+q5'length+q6'length downto 0+1+q1'length+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+1+q4'length downto 0+q0'length+q1'length+1+1);
q5 :=x(-1+q0'length+q1'length+1+1+q4'length+q5'length downto 0+q0'length+q1'length+1+1+q4'length);
q6 :=x(-1+q0'length+q1'length+1+1+q4'length+q5'length+q6'length downto 0+q0'length+q1'length+1+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+1+q4'length downto 0+1+1+q2'length+1);
q5 :=x(-1+1+1+q2'length+1+q4'length+q5'length downto 0+1+1+q2'length+1+q4'length);
q6 :=x(-1+1+1+q2'length+1+q4'length+q5'length+q6'length downto 0+1+1+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+1+q4'length downto 0+q0'length+1+q2'length+1);
q5 :=x(-1+q0'length+1+q2'length+1+q4'length+q5'length downto 0+q0'length+1+q2'length+1+q4'length);
q6 :=x(-1+q0'length+1+q2'length+1+q4'length+q5'length+q6'length downto 0+q0'length+1+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+1+q4'length downto 0+1+q1'length+q2'length+1);
q5 :=x(-1+1+q1'length+q2'length+1+q4'length+q5'length downto 0+1+q1'length+q2'length+1+q4'length);
q6 :=x(-1+1+q1'length+q2'length+1+q4'length+q5'length+q6'length downto 0+1+q1'length+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+1+q4'length downto 0+q0'length+q1'length+q2'length+1);
q5 :=x(-1+q0'length+q1'length+q2'length+1+q4'length+q5'length downto 0+q0'length+q1'length+q2'length+1+q4'length);
q6 :=x(-1+q0'length+q1'length+q2'length+1+q4'length+q5'length+q6'length downto 0+q0'length+q1'length+q2'length+1+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(0+1+1);
q3 :=x(-1+1+1+1+q3'length downto 0+1+1+1);
q4 :=x(-1+1+1+1+q3'length+q4'length downto 0+1+1+1+q3'length);
q5 :=x(-1+1+1+1+q3'length+q4'length+q5'length downto 0+1+1+1+q3'length+q4'length);
q6 :=x(-1+1+1+1+q3'length+q4'length+q5'length+q6'length downto 0+1+1+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(0+q0'length+1);
q3 :=x(-1+q0'length+1+1+q3'length downto 0+q0'length+1+1);
q4 :=x(-1+q0'length+1+1+q3'length+q4'length downto 0+q0'length+1+1+q3'length);
q5 :=x(-1+q0'length+1+1+q3'length+q4'length+q5'length downto 0+q0'length+1+1+q3'length+q4'length);
q6 :=x(-1+q0'length+1+1+q3'length+q4'length+q5'length+q6'length downto 0+q0'length+1+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(0+1+q1'length);
q3 :=x(-1+1+q1'length+1+q3'length downto 0+1+q1'length+1);
q4 :=x(-1+1+q1'length+1+q3'length+q4'length downto 0+1+q1'length+1+q3'length);
q5 :=x(-1+1+q1'length+1+q3'length+q4'length+q5'length downto 0+1+q1'length+1+q3'length+q4'length);
q6 :=x(-1+1+q1'length+1+q3'length+q4'length+q5'length+q6'length downto 0+1+q1'length+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+1+q3'length downto 0+q0'length+q1'length+1);
q4 :=x(-1+q0'length+q1'length+1+q3'length+q4'length downto 0+q0'length+q1'length+1+q3'length);
q5 :=x(-1+q0'length+q1'length+1+q3'length+q4'length+q5'length downto 0+q0'length+q1'length+1+q3'length+q4'length);
q6 :=x(-1+q0'length+q1'length+1+q3'length+q4'length+q5'length+q6'length downto 0+q0'length+q1'length+1+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(0+1);
q2 :=x(-1+1+1+q2'length downto 0+1+1);
q3 :=x(-1+1+1+q2'length+q3'length downto 0+1+1+q2'length);
q4 :=x(-1+1+1+q2'length+q3'length+q4'length downto 0+1+1+q2'length+q3'length);
q5 :=x(-1+1+1+q2'length+q3'length+q4'length+q5'length downto 0+1+1+q2'length+q3'length+q4'length);
q6 :=x(-1+1+1+q2'length+q3'length+q4'length+q5'length+q6'length downto 0+1+1+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(0+q0'length);
q2 :=x(-1+q0'length+1+q2'length downto 0+q0'length+1);
q3 :=x(-1+q0'length+1+q2'length+q3'length downto 0+q0'length+1+q2'length);
q4 :=x(-1+q0'length+1+q2'length+q3'length+q4'length downto 0+q0'length+1+q2'length+q3'length);
q5 :=x(-1+q0'length+1+q2'length+q3'length+q4'length+q5'length downto 0+q0'length+1+q2'length+q3'length+q4'length);
q6 :=x(-1+q0'length+1+q2'length+q3'length+q4'length+q5'length+q6'length downto 0+q0'length+1+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic) is
begin
q0 :=x(0);
q1 :=x(-1+1+q1'length downto 0+1);
q2 :=x(-1+1+q1'length+q2'length downto 0+1+q1'length);
q3 :=x(-1+1+q1'length+q2'length+q3'length downto 0+1+q1'length+q2'length);
q4 :=x(-1+1+q1'length+q2'length+q3'length+q4'length downto 0+1+q1'length+q2'length+q3'length);
q5 :=x(-1+1+q1'length+q2'length+q3'length+q4'length+q5'length downto 0+1+q1'length+q2'length+q3'length+q4'length);
q6 :=x(-1+1+q1'length+q2'length+q3'length+q4'length+q5'length+q6'length downto 0+1+q1'length+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

procedure f_unpack7 (
x: in std_logic_vector;
q6: out std_logic_vector;
q5: out std_logic_vector;
q4: out std_logic_vector;
q3: out std_logic_vector;
q2: out std_logic_vector;
q1: out std_logic_vector;
q0: out std_logic_vector) is
begin
q0 :=x(-1+q0'length downto 0);
q1 :=x(-1+q0'length+q1'length downto 0+q0'length);
q2 :=x(-1+q0'length+q1'length+q2'length downto 0+q0'length+q1'length);
q3 :=x(-1+q0'length+q1'length+q2'length+q3'length downto 0+q0'length+q1'length+q2'length);
q4 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length downto 0+q0'length+q1'length+q2'length+q3'length);
q5 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length+q5'length downto 0+q0'length+q1'length+q2'length+q3'length+q4'length);
q6 :=x(-1+q0'length+q1'length+q2'length+q3'length+q4'length+q5'length+q6'length downto 0+q0'length+q1'length+q2'length+q3'length+q4'length+q5'length);
end f_unpack7;

end pack_unpack_pkg;
